module and_test(input A, input B, output Result);
    assign Result = A & B; // Bitwise AND operation
endmodule